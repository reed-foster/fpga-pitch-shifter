// input_queue.v - Reed Foster
// overlapped window generator; feeds frames to FFT module

module input_queue
    ( // ports
        input clock, reset_n,
        input input_valid,
        input [11:0] data_in,
        output [20:0] data_out,
        output output_valid, output_last
    );
    // architecture

endmodule
