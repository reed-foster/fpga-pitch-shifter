// adc.v - Reed Foster
// xadc wrapper

module adc
    ( // ports
        input clock, reset_n,
        input vauxn3, vauxp3,
        output [11:0] sampled_data,
        output data_valid
    );
    // architecture

endmodule
